library verilog;
use verilog.vl_types.all;
entity media_movel2_vlg_vec_tst is
end media_movel2_vlg_vec_tst;
